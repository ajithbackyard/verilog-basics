module notgate(output wire Y,
                             input wire A);
              not(Y,A);
endmodule