module andgate(output wire Y,
                             input wire A,B);
              
endmodule
