module xorgate(output wire Y,
                             input wire A,B);
              
endmodule
