module orgate(output wire Y,
                             input wire A,B);
              or (Y,A,B);
endmodule

