module notgate(output wire Y,
                             input wire A);
              
endmodule
