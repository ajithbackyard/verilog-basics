module xorgate(output wire Y,
                             input wire A,B);
              xor (Y,A,B);
endmodule
