module orgate(output wire Y,
                             input wire A,B);
              
endmodule

