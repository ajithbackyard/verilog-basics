module andgate(output wire Y,
                             input wire A,B);
              and (Y,A,B);
endmodule